library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity audiomatrix_tb is
end entity audiomatrix_tb;

architecture test of audiomatrix_tb is
	constant CLOCK_PERIOD : time := 8064 ps;	-- 124 MHz clock

	component audiomatrix_ram_write is
		port (
			clk					: in std_logic;
			sync_in				: in std_logic;
			input_data			: in std_logic_vector(112 * 24 - 1 downto 0);
			
			o_ram_write_addr	: out unsigned(6 downto 0);
			o_ram_data			: out std_logic_vector(24 - 1 downto 0);
			o_ram_wr_en			: out std_logic;
			o_write_done		: out std_logic
		);
	end component;
	
	component audiomatrix_ram is
		port (
			clk					: in std_logic;
			read_addr			: in unsigned(6 downto 0);
			write_addr			: in unsigned(6 downto 0);
			i_data				: in std_logic_vector(24 - 1 downto 0);
			wr_en				: in std_logic;

			o_data				: out  std_logic_vector(24 - 1 downto 0)
		);
	end component;
  
	component audiomatrix_ram_read is
		port (
			clk					: in std_logic;
			sync_in				: in std_logic;
			select_lines		: in std_logic_vector(112 * 8 - 1 downto 0);
			i_ram_data			: in std_logic_vector(24 - 1 downto 0);
			
			o_ram_read_addr		: out unsigned(6 downto 0);
			output_data			: out std_logic_vector(112 * 24 - 1 downto 0)
		);
	end component;

	signal tb_clk				: std_logic := '0';
	signal tb_sync_in			: std_logic := '0';
	signal tb_input_data		: std_logic_vector(112 * 24 - 1 downto 0) := "101010101010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000";
	
	-- Testrounting:
	-- Ch1 <- Input 1 (23 downto 0)
	-- Ch2 <- Input 1 (47 downto 24)
	-- Ch3 <- Input 2 (71 downto 48)
	-- Ch 112 <- Input 112
	signal tb_select_lines		: std_logic_vector(112 * 8 - 1 downto 0) := "01101111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000";
	signal tb_i_ram_data		: std_logic_vector(24 - 1 downto 0) := (others => '0');
	signal tb_o_ram_read_addr	: unsigned(6 downto 0);
	signal tb_o_ram_write_addr	: unsigned(6 downto 0);
	signal tb_o_ram_data		: std_logic_vector(24 - 1 downto 0);
	signal tb_o_ram_wr_en		: std_logic;
	signal tb_o_write_done		: std_logic;
	signal tb_output_data		: std_logic_vector(112 * 24 - 1 downto 0);
begin
	-- Reset and clock
	tb_clk <= not tb_clk after CLOCK_PERIOD/2;
	tb_sync_in <= '0', '1' after (CLOCK_PERIOD/2), '0' after 2*(CLOCK_PERIOD/2), '1' after 5167*(CLOCK_PERIOD/2), '0' after 5169*(CLOCK_PERIOD/2), '1' after 10334*(CLOCK_PERIOD/2), '0' after 10336*(CLOCK_PERIOD/2);

--	tb_select_lines(tb_select_lines'high downto tb_select_lines'length - 8) <= std_logic_vector(to_unsigned(111, 8));
--	tb_select_lines(15 downto 8) <= std_logic_vector(to_unsigned(1, 8));

	-- declare the DUT modules
	dut1 : audiomatrix_ram_write
    port map (
		clk					=> tb_clk,
		sync_in				=> tb_sync_in,
		input_data			=> tb_input_data,

		o_ram_write_addr	=> tb_o_ram_write_addr,
		o_ram_data			=> tb_o_ram_data,
		o_ram_wr_en			=> tb_o_ram_wr_en,
		o_write_done		=> tb_o_write_done
    );
	
	dut2 : audiomatrix_ram
	port map (
		clk					=> tb_clk,
		read_addr			=> tb_o_ram_read_addr,
		write_addr			=> tb_o_ram_write_addr,
		i_data				=> tb_o_ram_data,
		wr_en				=> tb_o_ram_wr_en,

		o_data				=> tb_i_ram_data
	);

	dut3 : audiomatrix_ram_read
    port map (
		clk					=> tb_clk,
		sync_in				=> tb_o_write_done,
		select_lines		=> tb_select_lines,
		i_ram_data			=> tb_i_ram_data,

		o_ram_read_addr		=> tb_o_ram_read_addr,
		output_data			=> tb_output_data
    );
end architecture test;