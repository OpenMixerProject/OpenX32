`timescale 100 ps/100 ps
module ODDRX1F (
  SCLK,
  RST,
  D0,
  D1,
  Q
)
;
input SCLK ;
input RST ;
input D0 ;
input D1 ;
output Q ;
endmodule /* ODDRX1F */

